module counter_99 (count, clk, reset);
input clk;
input reset;
output reg [7:0] count;
endmodule